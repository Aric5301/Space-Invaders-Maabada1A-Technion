module	splashScreensBMP	(	
					input	logic	clk,
					input	logic	resetN,
					input logic	[10:0] offsetX,// offset from top left  position 
					input logic	[10:0] offsetY,
					input	logic	InsideRectangle, //input that the pixel is within a bracket 
					input logic [1:0] splashMode,

					output logic drawingRequest, //output that the pixel should be dispalyed 
					output logic [7:0] RGBout  //rgb value from the bitmap 
 );
 

// Size represented as Number of X and Y bits 
localparam logic [7:0] TRANSPARENT_ENCODING = 8'hFF ;// RGB value in the bitmap representing a transparent pixel 
 /*  end generated by the tool */


// the screen is 640*480  or  20 * 15 squares of 32*32  bits ,  we wiil round up to 32*16 and use only the top left 20*15 pixels  
// this is the bitmap  of the maze , if there is a one  the na whole 32*32 rectange will be drawn on the screen 
// all numbers here are hard coded to simplify the  understanding 
 
logic [0:2] [0:15] [0:127] [7:0] object_colors = {
{{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'h49,8'hFF,8'h49,8'h49,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'hFF,8'hFF,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h49,8'h49,8'h49,8'h49,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}
},
{{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hc0,8'hc0,8'hc0,8'hc0,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}
},
{{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'hFF,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'h18,8'h18,8'h18,8'h18,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF},
{8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF,8'hFF}
}};
 

// pipeline (ff) to get the pixel color from the array 	 

//==----------------------------------------------------------------------------------------------------------------=
always_ff@(posedge clk or negedge resetN) begin
	
	if(!resetN) begin
		RGBout <= 8'h00;
	end
	
	else begin
		RGBout <= TRANSPARENT_ENCODING ; // default 

		if ((InsideRectangle == 1'b1)) 
			RGBout <= object_colors[splashMode][offsetY][offsetX] ; 
		end 
end

//==----------------------------------------------------------------------------------------------------------------=
// decide if to draw the pixel or not 
assign drawingRequest = (RGBout != TRANSPARENT_ENCODING) ? 1'b1 : 1'b0 ; // get optional transparent command from the bitmpap   
endmodule